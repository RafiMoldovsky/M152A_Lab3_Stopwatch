`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:38:33 02/08/2022 
// Design Name: 
// Module Name:    stopwatch_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module stopwatch_tb();
//inputs 
reg clk;

//outputs
reg [7:0] seg;
reg [3:0] an;

stopwatch stopwatch_uut(.clk(clk),.seg(seg),.an(an));

initial begin
    clk=0;
    seg=8'b11111111;
    an=4'b1111;
end

always begin
    clk=~clk;
end

endmodule
